library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity DECODING_UNIT is
    port(
    DECODING_UNIT_in_INSTR    : in  std_logic_vector(31 downto 0));
end entity DECODING_UNIT;

architecture BEHAVIORAL of DECODING_UNIT is
    
begin

end architecture BEHAVIORAL;
