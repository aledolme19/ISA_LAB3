---------------------------------------------------------------------------------------------
-- File: IMM_UNIT.vhd
---------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity CONTROL_UNIT is
    port(
 
    );
end entity CONTROL_UNIT;

architecture BEHAVIORAL of CONTROL_UNIT is

begin



end BEHAVIORAL;