---------------------------------------------------------------------------------------------
-- File: IMM_UNIT.vhd
---------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity IMM_UNIT is
    port(
 
    );
end entity IMM_UNIT;

architecture BEHAVIORAL of IMM_UNIT is

begin



end BEHAVIORAL;