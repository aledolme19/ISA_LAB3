---------------------------------------------------------------------------------------------
-- File: RISC_V.vhd
---------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity RISC_V is
    port(
        clk : in std_logic
    );
end entity RISC_V;

architecture BEHAVIORAL of RISC_V is

begin

end BEHAVIORAL;
